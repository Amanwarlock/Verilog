

module Controller();

endmodule