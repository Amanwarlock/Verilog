module Multiplier256 #(
	parameter WIDTH = 256,
	parameter N = 2
)(
	input clk,
	input [WIDTH-1:0] a,b,
	output reg [2*WIDTH-1:0] prod
);

always @(clk) begin
	prod = a * b;
end



endmodule
