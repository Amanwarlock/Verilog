
module Gcd();

endmodule
